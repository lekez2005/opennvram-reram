.subckt sky130_fd_pr__reram_reram_cell TE BE
.param area_ox=0.1024e-12
Xreram TE BE state_out reram_cell_model area_ox='area_ox'
.ends
